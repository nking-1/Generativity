(** * Core Module - Re-exports all core DAO types
    
    This module provides a single import point for all the core types
    in the DAO framework: OmegaType, AlphaType, NomegaType, and GenerativeType.
*)

(** Re-export all core types *)
Require Export DAO.Core.OmegaType.
Require Export DAO.Core.AlphaType.
Require Export DAO.Core.NomegaType.
Require Export DAO.Core.GenerativeType.

(** ** The DAO Framework Summary
    
    - OmegaType: Complete but paradoxical (contains everything)
    - NomegaType: Empty but equally trivial (contains nothing) 
    - AlphaType: Consistent but incomplete (omega_veil maintains structure)
    - GenerativeType: Adds time dimension to resolve paradoxes temporally
    
    The omega_veil boundary prevents the collapse from Alpha to Omega/Nomega,
    maintaining the gradient that enables mathematics and meaning.
*)